-- PCS3412 - Organizacao e Arquitetura de Computadores I
-- PicoMIPS
-- File: ICache.vhd
-- Author: Daniel Nery Silva de Oliveira
--
-- Description:
--     Cache para Memoria de instrucoes

entity ICache is

end entity ICache;

architecture ICache_arch of ICache is

begin

end architecture ICache_arch;
