-- Testbench
-- Joins PC, ICache, MP and RI to test instruction fetch


entity instruction_fetch_tb is
end instruction_fetch_tb;

architecture instruction_arch of instruction_fetch_tb is

begin

end instruction_arch;
